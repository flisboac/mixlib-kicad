* ADA4522-4
* Packages: SOIC-14, TSSOP-14
* Pins:
*  1: OUT_A
*  2: -IN_A
*  3: +IN_A
*  4: V- (VIN-)
*  5: +IN_B
*  6: -IN_B
*  7: OUT_B
*  8: OUT_C
*  9: -IN_C
* 10: +IN_C
* 11: V+ (VIN+)
* 12: +IN_D
* 13: -IN_D
* 14: OUT_D
.SUBCKT ADA4522-4 OUTA INA- INA+ V- INB+ INB- OUTB OUTC INC- INC+ V+ IND+ IND- OUTD
.include ./include/ADA4522.cir
X1 INA+ INA- V+ V- OUTA ADA4522
X2 INB+ INB- V+ V- OUTB ADA4522
X3 INC+ INC- V+ V- OUTC ADA4522
X4 IND+ IND- V+ V- OUTD ADA4522
.ENDS ADA4522-4
