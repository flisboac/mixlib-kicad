* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*---------- DMC2990UDJQ Spice Model ----------

.SUBCKT DMC2990UDJQ S1 G1 D2 S2 G2 D1
M1 D1 G1 S1 DMC2990UDJQ_NMOS
M2 D2 G2 S2 DMC2990UDJQ_PMOS
.ENDS DMC2990UDJQ

*NMOS
.SUBCKT DMC2990UDJQ_NMOS 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3  NMOS  L = 1E-006  W = 1E-006 
RD 10 1 0.3743 
RS 30 3 0.001 
RG 20 2 113 
CGS 2 3 2.5E-011 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1  VFB 1 
CGD 13 14 8E-011 
R1 13 0 1 
D1 12 13  DLIM 
DDG 15 14  DCGD 
R2 12 15 1 
D2 15 0  DLIM 
DSD 3 10  DSUB 
.MODEL NMOS NMOS  LEVEL = 3  VMAX = 1E+006  ETA = 0.01  VTO = 0.8716 
+ TOX = 6E-008  NSUB = 1.886E+016  KP = 2.108  U0 = 400  KAPPA = 10.7 
.MODEL DCGD D  CJO = 1.594E-011  VJ = 0.2646  M = 0.429 
.MODEL DSUB D  IS = 2.265E-009  N = 1.422  RS = 1.834  BV = 25  CJO = 2.7E-012  VJ = 0.2048  M = 0.1841 
.MODEL DLIM D  IS = 0.0001 
.ENDS


*PMOS
.SUBCKT DMC2990UDJQ_PMOS 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 0.6562 
RS 30 3 0.001 
RG 20 2 400 
CGS 2 3 2.653E-011 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 5.8E-011 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 0.001 
+ TOX = 6E-008 NSUB = 1E+016 KP = 0.6965 KAPPA = 32.11 VTO = -0.6305 
.MODEL DCGD D CJO = 1.549E-011 VJ = 0.1652 M = 0.3749 
.MODEL DSUB D IS = 3.478E-007 N = 2.097 RS = 3.705 
+ BV = 25 CJO = 3.247E-012 VJ = 1.719E-014 M = 0.02141 
.MODEL DLIM D IS = 0.0001 
.ENDS

*Diodes DMC2990UDJQ Spice Model v1.0 Last Revised 2016/9/21
