* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*
*DIODES_INC_SPICE_MODEL
*ORIGIN=DZSL_DPG_GM
*SIMULATOR=PSPICE
*DATE=10FEB2011
*VERSION=1
*PIN_ORDER         
* 1=E1    6=C1
* 2=B1    5=B2
* 3=C2    4=E2
*
.SUBCKT MMDT5401 E1 B1 C2 E2 B2 C1
Q1 C1 B1 E1 Mod1
Q2 C2 B2 E2 Mod1
*
.MODEL Mod1 PNP IS=6E-14 NF=1 BF=130 VAF=360 ISE=6E-14
+ NE=1.5 NR=1 BR=6.5 VAR=37 ISC=8E-12 NC=1.35 RC=0.08 RB=1 RE=0.25
+ CJC=13E-12 MJC=0.46  VJC=0.7 CJE=63E-12 MJE=0.41 VJE=0.9 
+ TF=6.7E-10 TR=1.03E-6 XTB=1.5 QUASIMOD=1 RCO=14 GAMMA=1.5E-8
.ENDS MMDT5401
*
*$