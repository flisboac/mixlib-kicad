* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*
*DIODES_INC_SPICE_MODEL
*ORIGIN=DZSL_DPG_GM
*SIMULATOR=PSPICE
*DATE=23JUL2010
*VERSION=1
*PIN_ORDER         P1=C1, P2=B1, P3=C2, P4=E2, P5=B2, P6=E1
*
.SUBCKT ZXTD4591E6 C1 B1 C2 E2 B2 E1
Q1 C1 B1 E1 ZXTD4591E6_NPN
Q2 C2 B2 E2 ZXTD4591E6_PNP
.ENDS ZXTD4591E6

.MODEL ZXTD4591E6_NPN NPN IS=3.05E-13 NF=1.0034 BF=200 IKF=0.8 VAF=165
+ ISE=8.0191E-14 NE=1.4126 NR=1.001 BR=50 IKR=0.6 VAR=69
+ ISC=1.6E-12 NC=1.38 RB=0.065 RE=0.109 RC=0.075
+ CJC=17.2E-12 MJC=0.3429 VJC=0.4298 CJE=96E-12
+ TF=0.71E-9 TR=2.5E-9

.MODEL ZXTD4591E6_PNP PNP IS =3.2E-14 BF =170 VAF=45 NF =0.977 IKF=1.25 ISE=7E-15
+ NE =1.35 BR =50 VAR=50 NR =.986 IKR=0.15 ISC=0.9E-14 NC =1.08 RB =0.16
+ RE =0.195 RC =0.185 CJE=104E-12 TF =0.7E-9 CJC=30.5E-12 TR =3E-9 VJC=0.395
+ MJC=0.415
*
*$
