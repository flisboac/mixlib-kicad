* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.


.SUBCKT DMC62D2SV S1 G1 D2 S2 G2 D1
M1 D1 G1 S1 DMC62D2SV_NMOS
M2 D2 G2 S2 DMC62D2SV_PMOS
.ENDS DMC62D2SV

*---------- DMC62D2SV_NMOS Spice Model ----------
.SUBCKT DMC62D2SV_NMOS D=10 G=20 S=30 
* TERMINALS : D G S
* MODEL FORMAT : SPICE3
* Editor : Stan Li
M1 1 2 3 3 NMOS L = 1E-006 W = 1E-006 
RD 10 1 0.87 
RS 30 3 0.0001 
RG 20 2 146.4 
CGS 2 3 4.431E-011 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1 VFB 1 
CGD 13 14 8.535E-011 
R1 13 0 1 
D1 12 13 DLIM 
DDG 15 14 DCGD 
R2 12 15 1 
D2 15 0 DLIM 
DSD 3 10 DSUB 
DESD1 2 5 DESD 
DESD2 3 5 DESD 
.MODEL DESD D BV = 21 
.MODEL NMOS NMOS LEVEL = 3 VMAX = 1E+005 ETA = 0 VTO = 1.681 
+ TOX = 1E-007 NSUB = 9.974E+015 KP = 1.05 U0 = 100 KAPPA = 0.2 IS = 0 
.MODEL DCGD D CJO = 5.861E-012 VJ = 0.5 M = 0.3886 
.MODEL DSUB D IS = 3.5E-011 N = 1.333 RS = 0.1033 BV = 76.93 
+ CJO = 1.93E-011 VJ = 0.6 M = 0.4466 XTI = 0 TT = 9.215E-009 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes Spice Model v1.2 Last Revised 2023/03/08

*---------- DMC62D2SV_PMOS Spice Model ----------
.SUBCKT DMC62D2SV_PMOS D=10 G=20 S=30 
* TERMINALS : D G S
* MODEL FORMAT : SPICE3
* Editor : Stan Li
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 2.054 
RS 30 3 0.0001 
RG 20 2 234.9 
CGS 2 3 3.232E-011 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 7.54E-011 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 750 VMAX = 1E+005 ETA = 0 IS = 0 
+ TOX = 1E-007 NSUB = 1E+016 KP = 1 KAPPA = 0.2 VTO = -1.631 
.MODEL DCGD D CJO = 1.6E-011 VJ = 0.6 M = 0.468 
.MODEL DSUB D IS = 4.3E-010 N = 1.611 RS = 0.1045 BV = 76.39 
+ CJO = 9E-012 VJ = 0.7797 M = 0.3 XTI = 0 TT = 1.341E-008 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes Spice Model v1.2 Last Revised 2023/03/07

*The model is an approximation of the device, and it may not show the true device performance under all conditions.
*The model only guarantees the accuracy of the key parameters (Ron, VSD, IDSS, Ciss, Coss, Crss, and Trr) at 25 degC in the current data sheet.