* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*---------- DMP6023LFG Spice Model ----------
.SUBCKT DMP6023LFG 10 20 30 
* TERMINALS : D G S
* MODEL FORMAT : SPICE3
* Editor : J
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 0.01765 
RS 30 3 0.0005 
RG 20 2 4.99 
CGS 2 3 2.67E-009 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 1.99E-009 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 600 VMAX = 1E+005 ETA = 0 IS = 0 
+ TOX = 1E-007 NSUB = 1E+015 KP = 77 KAPPA = 0.2 VTO = -2.42 
.MODEL DCGD D CJO = 7.065E-010 VJ = 0.5048 M = 0.3861 
.MODEL DSUB D IS = 2.6E-009 N = 1.355 RS = 0.003114 BV = 66.8 
+ CJO = 2.986E-010 VJ = 0.7323 M = 0.5633 XTI = 0 TT = 9.9E-009 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes Spice Model v1.1 Last Revised 2021/12/22