* ADA4522-2
* Packages: SOIC-8, MSSOP-8
* Pins:
*  1: OUT_A
*  2: -IN_A
*  3: +IN_A
*  4: V- (VIN-)
*  5: +IN_B
*  6: -IN_B
*  7: OUT_B
*  8: V+ (VIN+)
.SUBCKT ADA4522-2 OUTA INA- INA+ V- INB+ INB- OUTB V+
.include ./include/ADA4522.cir
X1 INA+ INA- V+ V- OUTA ADA4522
X2 INB+ INB- V+ V- OUTB ADA4522
.ENDS ADA4522-2
