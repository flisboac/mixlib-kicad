* ADA4522-4 SPICE Macro-model
* Description: Amplifier
* Generic Desc: HV, ZD, Low Noise, Non-RRin, RRout
* Developed by: JG ADGT / VW ADSJ
* Revision History: 
* 05/18/2015 - initial release for dual
* 10/27/2015 - initial release for quad
* 9/6/2017 - added current noise block
* 0.0 (05/2015)
* 1.0 (09/2017)
* Copyright 2015 by Analog Devices
* T=25�C
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
*$
.SUBCKT ADA4522         1   2   99  50  45
*#ASSOC Category=Op-amp symbol=opamp
*
* INPUT STAGE
*
M1   4  7  8  8 PIX L=1E-6 W=1.18E-04
M2   6  2  8  8 PIX L=1E-6 W=1.18E-04
M3  14  7 18 18 NIX L=1E-6 W=1.18E-04
M4  16  2 18 18 NIX L=1E-6 W=1.18E-04
RD1  4 50 1.33E+04
RD2  6 50 1.33E+04
RD3 99 14 1.33E+04
RD4 99 16 1.33E+04
C1 4  6 6.7E-13
C2 14 16 6.7E-13
I1 99  8 3.00E-05
I2 18 50 3.00E-05
V1 99  9 2.113E+00 
V2 19 50 1.203E-01 
D1 8  9 DX
D2 19 18 DX
EOS 7 1 POLY(4) (73,98) (22,98) (81,98) (83,98) -9.1E-06 0.1 0.1 0.1 0.1
IOS 1  2 100E-12
V5 99 3 2.2
D5 1 3 DX
D6 50 1 DX
V6 99 100 2.2
D7 2 100 DX
D8 50 2 DX
Ccm1 1 50 35E-12
Ccm2 2 50 35E-12
Cdm 1 2 7.0E-12
*
*CMRR
*
E1  72 98 POLY(2) (1,98) (2,98) 0 5.25E-03 5.25E-03
R10 72 73 1.89E+02
R20 73 98 4.8E-01
C10 72 73 1.00E-06
*
* PSRR
*
EPSY 21 98 POLY(1) (99,50) -2.712E-00 2.4
RPS1 21 22 1.59E+05
RPS2 22 98 3.18E-01
CPS1 21 22 1.00E-06
*
*
* VOLTAGE NOISE REFERENCE
*
VN1 80 98 0
RN1 80 98  265E-05
HN  81 98 VN1 6.6E0
RNHH1 81 183 5.3
CHH1 183 98 1E-012
*
* CURRENT NOISE 
*
FIBIAS1 1 98 V21 800E-6 
V21 700 98 0
R28 700 98 .0167
D38 710 700 DIN
V22 710 98 0.2
FIBIAS2 2 98 V23 800E-6 
V23 720 98 0
R29 720 98 .0167
D39 730 720 DIN
V27 730 98 0.2
*
*BPF
*
EV5 83 98 VALUE = { V(203,98)+V(205,98) }
R94 204 98 300
L92 200 210 6.0e-006
C92 210 204 9e-011
R93 200 204 5.5E03 
EV4 205 98 204 98 10.5
EV3 203 98 202 98 5.5
R92 202 98 200    
L91 200 201 3.0e-005
C91 201 202 10e-010
R91 200 202 1E03
EV1 200 98 81 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) 805.1E-06 -1.55E-9
*
* GAIN STAGE
*
G1 98 30 POLY(2) (4,6) (14,16) 0 7.103E-03 7.103E-03
R1 30 98 1.00E+06
RZ 455 31 0.195E+00
CF 30 31 4.05E-9
EZ 455 98 (45,98) 1
V3 32 30 -7.5E-04
V4 30 33 -4.9E-04
D3 32 98 DX
D4 98 33 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=3E-6 W=20E-04
M6  45 47 50 50 NOX L=3E-6 W=40E-04
EG1 99 46 POLY(1) (98,30) 8.523E-01 1
EG2 47 50 POLY(1) (30,98) 8.523E-01 1
*EG1 99 46 POLY(1) (98,30) 8.523E-01 1
*EG2 47 50 POLY(1) (30,98) 8.523E-01 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=4.00E-05,VTO=-0.83,LAMBDA=0.047,RD=7)
.MODEL NOX NMOS (LEVEL=2,KP=4.00E-05,VTO=+0.83,LAMBDA=0.047,RD=38)
.MODEL PIX PMOS (LEVEL=2,KP=1.50E-05,VTO=-0.5,LAMBDA=0.047)
.MODEL NIX NMOS (LEVEL=2,KP=4.00E-05,VTO=0.5,LAMBDA=0.022)
.MODEL DX D(IS=1E-14,RS=0.1)
.MODEL DIN D(IS=1e-15,KF=3.18E-12)
*
*
.ENDS ADA4522

* ADA4522-1
* Packages: SOIC-8, MSSOP-8
* Pins:
*  1: N/C
*  2: -IN
*  3: +IN
*  4: V- (VIN-)
*  5: N/C
*  6: OUT
*  7: V+ (VIN+)
*  8: N/C
.SUBCKT ADA4522-1  2 3 4 6 7
X1 3 2 7 4 6 ADA4522
.ENDS ADA4522-1

* ADA4522-2
* Packages: SOIC-8, MSSOP-8
* Pins:
*  1: OUT_A
*  2: -IN_A
*  3: +IN_A
*  4: V- (VIN-)
*  5: _IN_B
*  6: -IN_B
*  7: OUT_B
*  8: V+ (VIN+)
.SUBCKT ADA4522-2 1 2 3 4 5 6 7 8
X1 3 2 8 4 1 ADA4522
X2 5 6 8 4 7 ADA4522
.ENDS ADA4522-2

* ADA4522-4
* Packages: SOIC-14, TSSOP-14
* Pins:
*  1: OUT_A
*  2: -IN_A
*  3: +IN_A
*  4: V- (VIN-)
*  5: +IN_B
*  6: -IN_B
*  7: OUT_B
*  8: OUT_C
*  9: -IN_C
* 10: +IN_C
* 11: V+ (VIN+)
* 12: +IN_D
* 13: -IN_D
* 14: OUT_D
.SUBCKT ADA4522-4 1 2 3 4 5 6 7 8 9 10 11 12 13 14
X1  3  2  4 11  1 ADA4522
X2  5  6  4 11  7 ADA4522
X3 10  9  4 11  8 ADA4522
X4 12 13  4 11 14 ADA4522
.ENDS ADA4522-4

*
*$
