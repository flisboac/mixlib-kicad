.SUBCKT AO3401A G S D
X1 D G S UNIT
.SUBCKT UNIT 4 1 2
M1  3 1 2 2 PMOS W=998956u  L=1.0u 
M2  2 1 2 4 NMOS W=998956u  L=0.7u
R1  4 3     RTEMP 17E-3
CGS 1 2     30E-12
DBD 3 2     DBD
**************************************************************************
.MODEL  PMOS       PMOS  (LEVEL  = 3               TOX    = 2.5E-8
+ RS     = 2E-4           RD     = 0               NSUB   = 2E17  
+ UO     = 120             THETA  = 0.2		   VTO=-1.1
+ VMAX   = 5e6             XJ     = 4E-7            KAPPA  = 1.2
+ ETA    = 0              TPG    = 1  
+ IS     = 0              LD     = 0                           
+ CGSO   = 0              CGDO   = 0               CGBO   = 0 
+ NFS    = 2E10         DELTA  = 0)
*************************************************************************
.MODEL  NMOS       NMOS (LEVEL   = 3               TOX    = 5.2E-8
+NSUB    = 2.0E16           TPG    = -1)   
*************************************************************************
.MODEL DBD D (CJO=900E-13     VJ=0.6    M=0.3
+RS=0.005 FC=0.5 IS=1E-12 TT=1.6E-8 N=1.0 BV=36 IBV=1E-4)
*************************************************************************
.MODEL RTEMP RES (TC1=1.5E-3   TC2=1E-6)
*************************************************************************
.ENDS UNIT
.ENDS AO3401A
