***********************************************************
*
* PBSS9110T
*
* Nexperia
*
* Low VCEsat PNP (BISS) Transistor
* IC   = 1 A
* VCEO = 100 V 
* hFE  = 150 - 450  @ 5V/500mA
*
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base
* Package Pin 2: Emitter
* Package Pin 3: Collector
*
*
* Extraction date (week/year): 31/2021
* Spicemodel includes temperature dependency
*
**********************************************************
*#
* Please note: Diode D1, Transistor Q2 and Resistor RQ 
* are dedicated to improve modeling of quasi
* saturation area and reverse mode operation
* and do not reflect physical devices.
*
.SUBCKT PBSS9110T B E C
Q1 B E C MAIN 0.8761
Q2 11 E C MAIN 0.1239
RQ B 11 26.15
D1 B E DIODE
*
.MODEL MAIN PNP
+ IS = 3.818E-13
+ NF = 0.9664
+ ISE = 5.361E-14
+ NE = 1.273
+ BF = 390.8
+ IKF = 0.8566
+ VAF = 40.32
+ NR = 0.9663
+ ISC = 1.16E-14
+ NC = 1.296
+ BR = 17.97
+ IKR = 8.103
+ VAR = 12.13
+ RB = 8
+ IRB = 0.001
+ RBM = 1.7
+ RE = 0.08877
+ RC = 0.03208
+ XTB = 0.5986
+ EG = 1.11
+ XTI = 1.368
+ CJE = 2.051E-10
+ VJE = 0.7516
+ MJE = 0.38
+ TF = 1.423E-09
+ XTF = 9.352
+ VTF = 1
+ ITF = 1.847
+ PTF = 0
+ CJC = 4.977E-11
+ VJC = 0.8642
+ MJC = 0.491
+ XCJC = 1
+ TR = 5.6E-08
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 1.288
.MODEL DIODE D
+ IS = 1.179E-13
+ N = 1.016
+ BV = 1000
+ IBV = 0.001
+ RS = 258.6
+ CJO = 0
+ VJ = 1
+ M = 0.9
+ FC = 0
+ TT = 0
+ EG = 1.1
+ XTI = 3
.ENDS PBSS9110T
*