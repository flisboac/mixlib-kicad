********************************
* Copyright:                   *
* Vishay Intertechnology, Inc. *
********************************
*Oct 09, 2017
*ECN S17-1578, Rev. A
*File Name: Si7223DN_PS.txt and Si7223DN_PS.lib
*This document is intended as a SPICE modeling guideline and does not
*constitute a commercial product datasheet. Designers should refer to the
*appropriate datasheet of the same number for guaranteed specification
*limits.
.SUBCKT SI7223DN S1 G1 S2 G2 D1 D2
X1 D1 G1 S1 Si7223DN
X2 D2 G2 S2 Si7223DN
.SUBCKT Si7223DN D G S 
M1 3 GX S S PMOS W= 2760000u L= 0.30u 
M2 S GX S D NMOS W= 2760000u L= 0.28u 
R1 D 3 1.840e-02 TC=3.985e-03,1.996e-06
CGS GX S 8.385e-10 
CGD GX D 8.387e-11 
RG G GY 8.6 
RTCV 100 S 1e6 TC=2.984e-03,3.034e-06
ETCV GY GX 100 200 1 
ITCV S 100 1u 
VTCV 200 S 1 
DBD D S DBD 2760000u 
*****************************************************  
.MODEL PMOS PMOS ( LEVEL = 3 TOX = 5e-8 
+ RS = 0 KP = 3.726e-06 NSUB = 3.304e+16 
+ KAPPA = 7.237e-03 NFS = 4.323e+11 
+ LD = 0 IS = 0 TPG = -1    )
***************************************************** 
.MODEL NMOS NMOS ( LEVEL = 3 TOX = 5e-8 
+NSUB = 1.963e+16 IS = 0 TPG = -1    )
***************************************************** 
.MODEL DBD D ( 
+FC = 0.1 TT = 1.001e-07 T_measured = 25 BV = 30.6
+RS = 2.919e-02 N = 1.096e+00 IS = 2.592e-12 
+EG = 8.778e-01 XTI = 9.824e+00 TRS1 = 3.133e-03
+CJO = 2.000e-11 VJ = 4.005e+00 M = 8.498e-01 ) 
.ENDS Si7223DN
.ENDS SI7223DN
