.SUBCKT MCP6407 VOUTA VINA- VINA+ VSS VINB+ VINB- VOUTB VDD
.include ./include/MCP640x.cir
X1 VINA+ VINA- VDD VSS VOUTA MCP640X
X2 VINB+ VINB- VDD VSS VOUTB MCP640X
.ENDS MCP6407
