.SUBCKT MCP6401R VOUT VDD VIN+ VIN- VSS
.include ./include/MCP640x.cir
X1 VIN+ VIN- VDD VSS VOUT MCP640X
.ENDS MCP6401R
