* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*ZETEX BSS138 Spice Model v2.0 Last Revised 5/4/07
*
.SUBCKT BSS138/ZTX D G S
* Nodes        D G S
M1 D 2 S S MOD1
RG G 2 20
RL D S 6E6
C1 2 S 30E-12
C2 D 2 1E-12 
C3 7 S 58E-12
D1 S D Dmod1
D2 6 D Dmod2
Egs1 2 6 2 S 1
Egs2 8 S 2 S 1
S1 2 7 D 2 SMOD1a
S2 7 8 D 2 SMOD1b
.MODEL MOD1 NMOS VTO=1 RS=1.58 RD=0.0 IS=1E-15 KP=0.395
+CBD=53.5E-12 PB=1 LAMBDA=267E-6
.MODEL Dmod1 D IS=1.254E-13 N=1.0207 RS=0.222
.MODEL Dmod2 D CJO=40E-12
.MODEL SMOD1a VSWITCH RON=1e-2 ROFF=1e4  VON=-1 VOFF=1
.MODEL SMOD1b VSWITCH RON=1e-2 ROFF=1e4  VON=1 VOFF=-1
.ENDS
*
*$
*

*BSS138 at Temp. Electrical Model
* Not ideal for Kicad
*-------------------------------------
* .SUBCKT BSS138 DRAIN GATE SOURCE VTEMP
* *20=DRAIN 10=GATE 30=SOURCE 50=VTEMP
* Rg GATE 11x 1
* Rdu 12x 1 1u
* M1 2 1 4x 4x DMOS L=1u W=1u
* .MODEL DMOS NMOS(VTO=1.35 KP=1.1
* +THETA=0.1 VMAX=1.5E5 LEVEL=3)
* Cgs 1 5x 22p
* Rd DRAIN 4 2.3E-1 
* Dds 5x 4 DDS
* .MODEL DDS D(M=3.93E-1 VJ=9.28E-1 CJO=29p)
* Dbody 5x DRAIN DBODY
* .MODEL DBODY D(IS=1.65E-10 N=1.413586 RS=.00148 TT=18.3n)
* Ra 4 2 2.3E-1
* Rs 5x 5 0.5m
* Ls 5 SOURCE 0.5n
* M2 1 8 6 6 INTER
* E2 8 6 4 1 2
* .MODEL INTER NMOS(VTO=0 KP=10 LEVEL=1)
* Cgdmax 7 4 118p
* Rcgd 7 4 10meg
* Dgd 6 4 DGD
* Rdgd 6 4 10meg
* .MODEL DGD D(M=5.05E-1 VJ=6.16E-2 CJO=118p)
* M3 7 9 1 1 INTER
* E3 9 1 4 1 -2
* *ZX SECTION
* EOUT 4x 6x poly(2) (1x,0) (3x,0) 0 0 0 0 1
* FCOPY 0 3x VSENSE 1
* RIN 1x 0 1G
* VSENSE 6x 5x 0
* RREF 3x 0 10m
* *TEMP SECTION
* ED 101 0 VALUE {V(50,100)}
* VAMB 100 0 25
* EKP 1x 0 101 0 .45
* *VTO TEMP SECTION
* EVTO 102 0 101 0 .001
* EVT 12x 11x 102 0 1
* *DIODE THEMO BREAKDOWN SECTION
* EBL VB1 VB2 101 0 .08
* VBLK VB2 0 VTEMP
* D DRAIN DB1 DBLK
* .MODEL DBLK D(IS=1E-14 CJO=.1p RS=.1)
* EDB DB1 0 VB1 0 1
* .ENDS BSS138
*BSS138 (Rev.A) 10/13/04 **ST


* NOTE: NOT supported in NGSPICE.
*
* BSS138 ELECTRICAL MODEL (SOT-23 Single N-Ch DMOS)
*-----------------------
* .SUBCKT  BSS138/FAI  20  10  30
* Rg     10    1    1
* M1      2    1    3    3    DMOS    L=1u   W=1u
* .MODEL DMOS NMOS (VTO={1.3*{-0.002*TEMP+1.05}}  KP={-0.0014*TEMP+0.685} THETA=0.086  VMAX=2.2E5  LEVEL=3)
* Cgs     1    3    40p
* Rd     20    4    0.2 TC=0.0065
* Dds     3    4    DDS
* .MODEL     DDS    D(BV={50*{0.00084*TEMP+0.979}}   M=0.36  CJO=23p   VJ=0.8)
* Dbody   3   20    DBODY
* .MODEL   DBODY    D(IS=1.4E-13   N=1   RS=40m   TT=100n)
* Ra      4    2    0.3 TC=0.0065
* Rs      3    5    10m
* Ls      5    30   .5n
* M2      1    8    6    6   INTER
* E2      8    6    4    1   2
* .MODEL   INTER    NMOS(VTO=0  KP=10   LEVEL=1)
* Cgdmax  7    4    68p
* Rcgd    7    4    10meg
* Dgd     6    4    DGD
* Rdgd    4    6    10meg
* .MODEL     DGD    D(M=0.3   CJO=68p   VJ=0.4)
* M3      7    9    1    1   INTER
* E3      9    1    4    1   -2
* .ENDS BSS138/FAI
