.SUBCKT MCP6406 VOUT VSS VIN+ VIN- VDD
.include ./include/MCP640x.cir
X1 VIN+ VIN- VDD VSS VOUT MCP640X
.ENDS MCP6406
