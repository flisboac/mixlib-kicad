.SUBCKT LM2903B 1OUT 1IN- 1IN+ GND 2IN+ 2IN- 2OUT V+
.include ./include/LM2903B.cir
X1 1IN+ 1IN- VCC GND 1OUT LM2903B
X2 2IN+ 2IN- VCC GND 2OUT LM2903B
.ENDS LM2903B
