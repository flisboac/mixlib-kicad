.SUBCKT LM4040_33  V+ V- PARAMS: TOL=0
C_Cstart         V- START  80nF  TC=0,0 
X_Q22        N06562 N10050 V- NPN1X PARAMS: AREA=1          
X_Q7         N06041 N05858 N06045 NPN1X PARAMS: AREA=1      
X_Q12         N06650 N06562 N06698 NPN1X PARAMS: AREA=1     
X_Q13         N06802 N06802 N06698 NPN1X PARAMS: AREA=10
X_Q3         N05681 VB_Q3 N05862 NPN1X PARAMS: AREA=10           
X_Q5         N05681 N06002 N01136 PNPL1X PARAMS: AREA = 1.34    
X_Q6         N06002 N06002 N01136 PNPL1X PARAMS: AREA = 1.8      
C_C3         N06562 N01136  3pF  TC=0,0    
X_Q23         N01136 N01136 N07802 NPN1X PARAMS: AREA=1
R_R10         N06002 N06045  60K TC=0,0    
X_Q15         N06802 N06650 N01136 PNPL1X PARAMS: AREA = 10      
R_R1toR5         N05442 N01136  30.5K TC=0,0            
R_R15         N10050 Q20B  66K TC=0,0     
X_Q14         N06650 N06650 N01136 PNPL1X PARAMS: AREA = 1      
X_Q20         N07708 Q20B V- NPN1X PARAMS: AREA=1
R_R6         VB_Q2 N05442  20K TC=0,0   
C_Cx         V- N01136  1pF  TC=0,0   
C_C2         N05681 N06272  6pF  TC=0,0   
X_Estart         N30465 V- VB_Q2  VB_Q3 Q20B  Estart   
X_Q1         V- N05136 N05430 PNPV1X PARAMS: AREA=5 
X_Q17         N07708 N05136 N05430 PNPL1X PARAMS: AREA = 1   
R_Rx6         N01137  N01136  500 TC=0,0 
R_R22         VX  N01137  0.100
R_R23         VX  N01147  0.096
L_Lx2         N01147  N01137 1000U
X_Q19         Q20B N05862 N08426 PNPL1X PARAMS: AREA = 1    
R_R8         N05430 VB_Q3  45K TC=0,0  
X_Q16         N01136 N06802 V- NPN1X PARAMS: AREA = 10   
X_Q4         N05858 N06002 N01136 PNPL1X PARAMS: AREA = 1.34
R_R13         Q20B N07708  40K TC=0,0     
R_Rstart0         START N30465  100 TC=0,0   
R_R11         N06272 N06041  100K TC=0,0     
R_R14         N06127 V-  3.3K TC=0,0         
X_Q11         N06562 N06272 N01136 PNPL1X PARAMS: AREA = 1.8   
X_Q21         N06045 Q20B N06127 NPN1X PARAMS: AREA=6.75  
X_Q24         N01136 N05442 N07806 NPN1X PARAMS: AREA=1    
X_Q8         N06272 N05681 N06045 NPN1X PARAMS: AREA=1       
X_Q2         N05858 VB_Q2 N05862 NPN1X             
X_Q10         N06272 N06041 N01136 PNPL1X PARAMS: AREA = 3.1
X_Q9         N06041 N06041 N01136 PNPL1X PARAMS: AREA = 3.1
R_R18         N05430 N07806  69K TC=0,0      
R_R59         N01136 N08426  51K TC=0,0   
R_R12         N05655 V-  6K TC=0,0    
L_Lx1         N01137 N01136  2.0uH  
R_R16         N06698 V-  1K TC=0,0      
X_Q18         N05862 Q20B N05655 NPN1X PARAMS: AREA=1
R_Rstart1         Q20B START  20K TC=0,0   
R_R17         N07806 N07802  130k TC=0,0 
R_R7         VB_Q3 VB_Q2  10K TC=0,0   
C_C1         N05858 N06562  3pF  TC=0,0    
X_R19       VX N05136  R_TOL PARAMS: RTOL = {TOL}   
R_R20       N05136 V-  800K     
X_U24       V+ VX V- VX  VCCS1       
R61     V+ VX 0.001

.subckt NPN1X 1 2 3  PARAMS: AREA = 1
Q1  1 2 3 _NPN1X {AREA}
.model _NPN1X	NPN Is=13.84e-18 Bf=130 TR=8ns
.ends NPN1X

.subckt PNPV1X 1 2 3  PARAMS: AREA = 1
Q1  1 2 3 _PNPV1X {AREA}
.model _PNPV1X	PNP Is=261.8e-18 Bf=222
.ends PNPV1X

.subckt PNPL1X 1 2 3  PARAMS: AREA = 1
Q1  1 2 3 _PNPL1X {AREA}
.model _PNPL1X	PNP  Is=48e-18 Bf=200
.ends PNPL1X

.subckt Estart 1 2 3 4 5
E_Estart    1 2 VALUE {max(0.4*(1-V(3, 4)/.05), 0)+V(5)}
.ends Estart

.subckt R_TOL 1 2 PARAMS: RTOL = 0
R_R1       1 2    {IF({RTOL}==0,469.42K,IF({RTOL}>0,467.94K,470.920K))}
.ends R_TOL

.SUBCKT VCCS1   VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {(V(VC+,VC-))} =
+(0,0u)
+(45n,-30u)
+(46n,0u)
+(47n,70u)
+(15u,70u)
.ENDS VCCS1

.ENDS  LM4040_33
*$
