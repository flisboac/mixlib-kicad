* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*****************************************************************************************************************************************
*SRC=MMDT4413;DI_MMDT4413_NPN;BJTs NPN; Si;  40.0V  0.600A  275MHz   Diodes Inc. BJTs - Complementaryl
.SUBCKT MMDT4413 E1 B1 C2 E2 B2 C1
X1 C1 B1 E1 MMDT4413_NPN
X2 C2 B2 E2 MMDT4413_PNP
.ENDS MMDT4413

.MODEL MMDT4413_NPN  NPN (IS=60.7f NF=1.00 BF=410 VAF=114
+ IKF=0.219 ISE=19.7p NE=2.00 BR=4.00 NR=1.00
+ VAR=24.0 IKR=0.540 RE=85.8m RB=0.343 RC=34.3m
+ XTB=1.5 CJE=36.2p VJE=1.10 MJE=0.500 CJC=15.4p VJC=0.300
+ MJC=0.300 TF=539p TR=84.1n EG=1.12 )

*SRC=MMDT4413;DI_MMDT4413_PNP;BJTs PNP; Si;  40.0V  0.600A  275MHz   Diodes Inc. BJTs - Complementary
.MODEL MMDT4413_PNP  PNP (IS=61.0f NF=1.00 BF=410 VAF=114
+ IKF=0.340 ISE=24.7p NE=2.00 BR=4.00 NR=1.00
+ VAR=20.0 IKR=0.840 RE=0.269 RB=1.08 RC=0.108
+ XTB=1.5 CJE=27.6p VJE=1.10 MJE=0.500 CJC=18.5p VJC=0.300
+ MJC=0.300 TF=516p TR=84.1n EG=1.12 )
*****************************************************************************************************************************************
