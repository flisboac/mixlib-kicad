***********************************************************
*
* PBSS8110T
*
* Nexperia
*
* Low VCEsat NPN (BISS) Transistor
* IC   = 1 A
* VCEO = 100 V 
* hFE  = 150 - 500  @ 10V/250mA
*
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base 
* Package Pin 2: Emitter
* Package Pin 3: collector
*
*
* Extraction date (week/year): 08/2004
* Spicemodel does not include temperature dependency
*
**********************************************************
*#
* Please note: Diode D1 is dedicated to improve modeling in reverse
* mode of operation and does not reflect a physical device.
*
.SUBCKT PBSS8110T B E C
Q1 B E C PBSS8110T
D1 E B DIODE
* 
.MODEL PBSS8110T NPN 
+ IS = 3.138E-013 
+ NF = 0.9857 
+ ISE = 4.405E-015 
+ NE = 1.299 
+ BF = 300 
+ IKF = 0.38 
+ VAF = 23 
+ NR = 0.9809 
+ ISC = 1.35E-016 
+ NC = 0.998 
+ BR = 55 
+ IKR = 2.8 
+ VAR = 48 
+ RB = 10 
+ IRB = 0.000431 
+ RBM = 5.92 
+ RE = 0.05 
+ RC = 0.058 
+ XTB = 0 
+ EG = 1.11 
+ XTI = 3 
+ CJE = 2.86E-010 
+ VJE = 0.7299 
+ MJE = 0.3486 
+ TF = 6E-010 
+ XTF = 27 
+ VTF = 1.5 
+ ITF = 0.6 
+ PTF = 0 
+ CJC = 2.39E-011 
+ VJC = 0.2734 
+ MJC = 0.3734 
+ XCJC = 1 
+ TR = 5.1E-008 
+ CJS = 0 
+ VJS = 0.75 
+ MJS = 0.333 
+ FC = 0.78 
.MODEL DIODE D 
+ IS = 1.185E-013 
+ N = 1 
+ BV = 1000 
+ IBV = 0.001 
+ RS = 500 
+ CJO = 0 
+ VJ = 1 
+ M = 0.5 
+ FC = 0 
+ TT = 0 
+ EG = 1.11 
+ XTI = 3 
.ENDS PBSS8110T
*