*Aug 13, 2012
*ECN S12-1928, Rev. A
*File Name: SUD50P06-15_PS.txt and SUD50P06-15_PS.lib
*This document is intended as a SPICE modeling guideline and does not
*constitute a commercial product datasheet. Designers should refer to the
*appropriate datasheet of the same number for guaranteed specification
*limits.
.SUBCKT SUD50P06-15 G D S
M1  3  G S S PMOS W=8943624u L=0.25u         
M2  S  G S D NMOS W=8943624u L=0.45u 
R1  D  3     RTEMP 5E-3
CGS G  S     3400E-12
DBD D  S     DBD
***************************************************************  
.MODEL  PMOS       PMOS  ( LEVEL  = 3           TOX    = 5E-8
+ RS     = 6.2E-3          RD     = 0           NSUB   = 1.05E17
+ KP     = 4E-6            UO     = 400             
+ VMAX   = 0               XJ     = 5E-7        KAPPA  = 5E-2
+ ETA    = 1E-4            TPG    = -1  
+ IS     = 0               LD     = 0                        
+ CGSO   = 0               CGDO   = 0           CGBO   = 0 
+ NFS    = 0.8E12          DELTA  = 0.1)
*************************************************************** 
.MODEL  NMOS       NMOS  ( LEVEL  = 3           TOX    = 5E-8
+NSUB    = 4E16            NFS    = 1E12        TPG    = -1)   
*************************************************************** 
.MODEL DBD D (CJO=200E-12 VJ=0.38 M=0.37
+RS=0.1 FC=0.5 IS=1E-12 TT=6E-8 N=1 BV=60.2)
*************************************************************** 
.MODEL RTEMP RES (TC1=13E-3 TC2=5.5E-6)
*************************************************************** 
.ENDS
