*******************************************************
* Taiwan Semiconductor
* SS16
* 1A, 60V Schottky Barrier Rectifier
* Date: 2023-05-04
*******************************************************
.SUBCKT SS16 K A
D1 A K SS16
.MODEL SS16 D
+ IS=57.136E-6
+ N=1.8535
+ RS=50.858E-3
+ IKF=.29449
+ CJO=126.83E-12
+ M=.51467
+ VJ=.52466
+ ISR=10.010E-21
+ NR=4.9950
+ BV=60
+ IBV=2E-4
+ TT=15.291E-9
.ENDS SS16
*******************************************************
