.SUBCKT LM358B-8PIN OUT1 IN1- IN1+ V- IN2+ IN2- OUT2 V+
.include ./include/LMx58B_LM2904B.cir
X1 IN1+ IN1- V+ V- OUT1 LMX58B_LM2904B
X2 IN2+ IN2- V+ V- OUT2 LMX58B_LM2904B
.ENDS LM358B-8PIN
