***********************************************************
*
* PBSS4160DS
*
* Nexperia
*
* Low VCEsat double NPN/NPN (BISS) Transistor
* Ic   = 1 A
* Vceo = 60 V 
* hFE  = min. 250 typ.500  @ 5V/1mA 
* 
*
* 
*
* Package pinning does not match Spice model pinning.
* Package: SOT 457
*  
* Package Pin 1;4: Emitter   TR1;TR2
* Package Pin 2;5: Base      TR1;TR2
* Package Pin 3;6: Collector TR2;TR1
*
*
* Extraction date (week/year): 31/2019
* Spicemodel includes temperature dependency
*
**********************************************************
*#
* Please note: The following model is to be used twice in 
* schematic due to equality of both Transistors.
*
* Diode D1 is dedicated to improve modeling in reverse
* mode of operation and does not reflect a physical device.
*
.SUBCKT PBSS4160DS E1 B1 C2 E2 B2 C1
X1 C1 B1 E1 PBSS4160DS_UNIT
X2 C1 B2 E2 PBSS4160DS_UNIT
.ENDS PBSS4160DS

.SUBCKT PBSS4160DS_UNIT 1 2 3
Q1 1 2 3 MAIN 
D1 2 1 DIODE 
*
.MODEL MAIN NPN 
+ IS = 1.903E-13
+ NF = 0.9792
+ ISE = 9.036E-16
+ NE = 1.126
+ BF = 503
+ IKF = 0.1644
+ VAF = 10
+ NR = 0.9805
+ ISC = 1E-18
+ NC = 1.821
+ BR = 50
+ IKR = 5.754
+ VAR = 18
+ RB = 19
+ IRB = 0.00043
+ RBM = 1.7
+ RE = 0.1259
+ RC = 0.1052
+ XTB = 0.9903
+ EG = 1.11
+ XTI = 0.7331
+ CJE = 1.115E-10
+ VJE = 0.587
+ MJE = 0.308
+ TF = 4.8E-10
+ XTF = 8
+ VTF = 1.5
+ ITF = 1.3
+ PTF = 0
+ CJC = 1.893E-11
+ VJC = 0.6185
+ MJC = 0.4452
+ XCJC = 1
+ TR = 4.3E-08
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 0.9
.MODEL DIODE D
+ IS = 8E-15
+ N = 0.98
+ BV = 1000
+ IBV = 0.001
+ RS = 850
+ CJO = 0
+ VJ = 1
+ M = 0.7
+ FC = 0
+ TT = 0
+ EG = 1.11
+ XTI = 3 
.ENDS PBSS4160DS_UNIT
*