* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*---------- DMG1029SV Spice Model ----------

.SUBCKT DMG1029SV S1 G1 D2 S2 G2 D1
M1 D1 G1 S1 DMG1029SV_N
M2 D2 G2 S2 DMG1029SV_P
.ENDS DMG1029SV

*NMOS
.SUBCKT DMG1029SV_N 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3  NMOS  L = 1E-006  W = 1E-006 
RD 10 1 1.631 
RS 30 3 0.001 
RG 20 2 133 
CGS 2 3 2.711E-011 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1  VFB 1 
CGD 13 14 2.628E-011 
R1 13 0 1 
D1 12 13  DLIM 
DDG 15 14  DCGD 
R2 12 15 1 
D2 15 0  DLIM 
DSD 3 10  DSUB 
.MODEL NMOS NMOS  LEVEL = 3  VMAX = 1E+006  ETA = 0  VTO = 1.596 
+ TOX = 6E-008  NSUB = 1.945E+017  KP = 1.196  KAPPA = 1E-015  U0 = 400  THETA = 5.648E-007 
.MODEL DCGD D  CJO = 2.628E-011  VJ = 0.009081  M = 0.2561 
.MODEL DSUB D  IS = 2.05E-009  N = 1.698  RS = 0.1282  BV = 65  CJO = 6.226E-012  VJ = 1  M = 0.6474 
.MODEL DLIM D  IS = 0.0001 
.ENDS

*PMOS
.SUBCKT DMG1029SV_P 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 2.072 
RS 30 3 0.001 
RG 20 2 50 
CGS 2 3 2.301E-011 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 4.1E-011 
R1 13 30 1 
D1 13 12  DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 0.001 TOX = 6E-008 NSUB = 1E+016 KP = 0.3083 KAPPA = 32.1 VTO = -1.513 
.MODEL DCGD D CJO = 7.698E-012 VJ = 0.2 M = 0.2205 
.MODEL DSUB D IS = 9.579E-010 N = 1.677 RS = 0.1623  BV = 65 CJO = 9.694E-012 VJ = 0.4761 M = 0.3849 
.MODEL DLIM D IS = 0.0001 
.ENDS

*Diodes DMG1029SV Spice Model v1.0 Last Revised 2012/4/17