.SUBCKT MCP6404 VOUTA VINA- VINA+ VDD VINB+ VINB- VOUTB VOUTC VINC- VINC+ VSS VIND+ VIND- VOUTD
.include ./include/MCP640x.cir
X1 VINA+ VINA- VDD VSS VOUTA MCP640X
X2 VINB+ VINB- VDD VSS VOUTB MCP640X
X3 VINC+ VINC- VDD VSS VOUTC MCP640X
X4 VIND+ VIND- VDD VSS VOUTD MCP640X
.ENDS MCP6404
