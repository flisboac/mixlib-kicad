* SPICE model Zener diodes ***ZMM1***
* Use the symbol file ***zmm1.asy***
*
* (c) Diotec Semiconductor AG
* www.diotec.com
* 2022-01-26
*
*********************************************************
* This model is for simulation purposes only. It does   *
* not replace reviewing of the data sheet nor real life *
* testing of the part inside the application.           *
*********************************************************
*
.subckt ZMMx  A  K  params: Vznom=0.765 Iztest=5m Vr=0.6 Ir=100u Rzj=8 Izmax=400m Cjo=700p

* Above values are an example for the ***ZMM1***. Using the
* above symbol file allows for direct insertion of other values
* according to these data sheet parameters:
*
* Vznom		Nominal zener voltage at 25�C = (Vzmin+Vzmax)/2
* Iztest	Test current for Vz
* Vr		Reverse voltage (minimum value)
* Ir		Reverse current
* Rzj		Dynamic resistance
* Izmax		Max zener current
* Cjo		Junction capacitance at 0V

Dbr  INT  K  Zbr
Df   A    K  Zf
Dbl  INT  A  DIObl

* Zener breakdown characteristic
.model  Zbr  D(Is={Ir/10} N=2.0 Rs={Rzj} Bv={Vznom*(1+(temp-25)*0.001)} Ibv={Iztest} Eg=1.11 Xti=3 M=.33 diss={Vznom*Izmax})
*
* Forward characteristic
.model  Zf  D(Is=100E-9 N=2.0 Rs=37m Cjo={Cjo} Eg=1.11 Xti=3 M=.33 Tt=800n)
*
* Internal blocking diode
.model  DIObl  D(Ron=.1m)

.ends ZMMx
