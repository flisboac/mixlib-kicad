.SUBCKT MCP6401U VIN+ VSS VIN- VOUT VDD
.include ./include/MCP640x.cir
X1 VIN+ VIN- VDD VSS VOUT MCP640X
.ENDS MCP6401U
