* source TPS61023
.SUBCKT TPS61023_Symbol FB EN VIN GND SW VOUT  
X_U1 EN FB GND SW VIN VOUT TPS61023_schematic  
.ENDS
 
.SUBCKT TPS61023_schematic EN FB GND SW VIN VOUT  
D_D5         VOUT_INT N03750 D_D1 
E_E1         N04714 0 VOUT_INT 0 0.3
R_R9         N03512 PRECHARGE_ON  1 TC=0,0 
X_S4    PRECHARGE_ON 0 SW N03792 TPS61023_schematic_S4 
X_H2    N03792 N03994 ISEN_LDO 0 TPS61023_schematic_H2 
X_S2    SDWN 0 N03792 N04226 TPS61023_schematic_S2 
X_U5 EN SDWN VIN VOUT Enable_UVLO  
D_D7         VOUT N03750 D_D1 
C_C10         N03994 N04226  208p IC={{SS}*2} TC=0,0 
D_D6         N04164 VOUT_INT D_D1 
X_S1    GATE_NMOS 0 SW 0 TPS61023_schematic_S1 
X_D1         0 SW D_Dnew 
V_V5         N04404 0 5
X_U2 GATE_NMOS GATE_PMOS OVP PASS_THROUGH PRECHARGE N02524 N02652 SDWN
+  SKIP_PFM_N Gate_Driver  
M_M1         VOUT_INT N04226 N03994 N03994 MbreakP           
G_ABM2I5         N04226 0 VALUE { {LIMIT((V(N04226) - V(VIN))*500u, 0,30u)}   
+  }
X_U1 FB_INT ISEN_LDO PFM PRECHARGE_ON VREF SDWN VEA Error_Amp  
E_ABM10         MAX 0 VALUE { max(V(VIN), V(VOUT))    }
X_F1    N02802 N02682 0 VOUT_INT TPS61023_schematic_F1 
X_U10         SDWN N03284 INV_BASIC_GEN PARAMS: VDD=1 VSS=0 VTHRESH=500E-3
G_ABM2I6         0 N04226 VALUE { {LIMIT((V(0) - V(N04226))*500u, 0,30u)}    }
X_U4 FB_INT PRECHARGE_ON SDWN VREF Soft_Start  
R_R8         N03590 PRECHARGE  1 TC=0,0 
X_U7 OVP VOUT OVP  
E_ABM176         N03428 0 VALUE { (V(VIN) -  200m)     }
X_U616         N03428 VOUT N03668 N03590 COMPHYS_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=0.5
D_D8         N04164 VOUT D_D1 
R_R7         0 N04226  200MEG TC=0,0 
V_V16         N02676 MAX 0.6
X_H1    SW N02802 ISENSE 0 TPS61023_schematic_H1 
X_U6 FB_INT PASS_THROUGH PRECHARGE_ON VIN VOUT Pass_Through  
G_ABM2I4         N04404 N04226 VALUE { {LIMIT((V(ISEN_LDO)*2 -
+  V(VOUT_SEN))*10u, -3u,3u)}    }
E_ABM174         VOUT_SEN 0 VALUE {  IF(V(N04714) > 180m, V(N04714),180m)    }
X_U11         N03284 PRECHARGE N03512 AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U9 FB_INT GATE_NMOS GATE_PMOS 0 PFM VREF SKIP_PFM SKIP_PFM_N VEA MODE_SKIP  
E_E2         FB_INT 0 N18081 0 1
D_D4         N02682 N02676 D_D1 
X_S3    GATE_PMOS 0 N02802 VOUT_INT TPS61023_schematic_S3 
C_C11         0 PRECHARGE  1n  TC=0,0 
X_U3 ISENSE GATE_PMOS N02524 N02652 SKIP_PFM VEA VIN VOUT PWM_Control  
I_I1         N03750 N04164 DC 10A  
C_C12         0 PRECHARGE_ON  5n  TC=0,0 
V_V17         N03668 0 2m
R_R10         FB N18081  50k TC=0,0 
C_C14         0 N18081  800f  TC=0,0 
C_C13         0 FB  1p  TC=0,0 
.ENDS
 
.SUBCKT PWM_Control ISENSE pMOS_GATE PWM PWM_N SKIP_PFM VEA VIN VOUT  
X_U22         N16760623 RESET PWM PWM_N SRLATCHRHP_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
E_ABM175         ISEN_INT 0 VALUE {  IF((V(N16805500) > 0.5) , V(ISENSE) ,   
+ 0)   }
C_C14         RESET 0  1n  TC=0,0 
X_U620         N16794413 TON_EXP RESET_INT AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U621         N16799638 N16798891 INV_DELAY_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=0.5 DELAY=10n
D_D2         N16760219 N16760209 D_D1 
R_R11         RESET_INT RESET  1 TC=0,0 
X_U624         PWM SKIP_N N16852133 AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
C_C13         N16788226 0  1.443n  TC=0,0 
X_U10 TON VIN VOUT ON_TIME_VALUE  
X_U625         PMOS_GATE BLNK_TIME N16805500 AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
C_C2         N16760219 0  1u  
X_U622         N16798891 N16799638 N16788246 AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
D_D4         BLNK_TIME PMOS_GATE D_D1 
X_U615         VEA ISEN_INT N167609210 N16760623 COMPHYS_BASIC_GEN PARAMS:
+  VDD=1 VSS=0 VTHRESH=0.5
E_E1         N16760203 0 TON 0 1000
X_U630         RESET_INT N16833195 ONE_SHOT PARAMS:  T=90  
X_U631         SKIP_PFM PWM_N N16851858 OR2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
G_ABMII1         N16760209 N16760219 VALUE { (V(N16852133) *1m)    }
D_D5         N16788246 N16788226 D_D1 
V_V7         N167609210 0 2m
V_V2         N16760209 0 2
X_U619         N16788226 N16794413 INV_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U629         N16760219 N16760203 N16834033 COMP_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=0.5
C_C12         BLNK_TIME 0  1.443n  TC=0,0 
X_U628         N16834033 N16833195 TON_EXP OR2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U626         PWM SKIP_N N16799638 AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U623         SKIP_PFM SKIP_N INV_BASIC_GEN PARAMS: VDD=1 VSS=0 VTHRESH=500E-3
X_S2    N16851858 0 N16760219 0 PWM_Control_S2 
R_R10         N16788246 N16788226  70 TC=0,0 
R_R9         PMOS_GATE BLNK_TIME  70 TC=0,0 
.ENDS
 
.SUBCKT ON_TIME_VALUE TON VIN VOUT  
E_ABM4         N00593 0 VALUE { TANH((V(VIN) -1.3)* 6.5)    }
E_ABM7         N01724 0 VALUE { (V(VOUT_P) *12000*3/(2*0.658e6))    }
E_ABM5         N00775 0 VALUE { (((V(N00593) +1)*0.5)+1)*0.5    }
E_ABM9         N03521 0 VALUE { (( V(N01998)  
+ / V(N00775) )+40n)   }
E_ABM6         VOUT_P 0 VALUE { (V(VOUT) +0.1)    }
E_ABM3         N00363 0 VALUE { ( V(VOUT)  
+ - V(VIN) )   }
C_C12         0 TON  1n  TC=0,0 
R_R9         N03521 TON  1 TC=0,0 
E_ABM8         N01998 0 VALUE { (( V(N00363)  
+ - V(N01724) )*1.974e-6/(2*V(VOUT_P)))   }
.ENDS
 
.SUBCKT MODE_SKIP FB_INT GATE_nMOS GATE_pMOS MODE PFM REF SKIP_PFM SKIP_PFM_N
+  VEA  
X_U623         SKIP PFM SKIP_PFM AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U628         N16788254 N16764440 N16786337 SKIP AND3_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=500E-3
X_U617         FPWM PFM INV_BASIC_GEN PARAMS: VDD=1 VSS=0 VTHRESH=500E-3
C_C1         N16761926 0  1p  TC=0,0 
E_E1         N16761940 0 REF 0 1.01
V_V6         N16763091 0 50u
X_U619         N16763641 VEA N16763659 N16764440 COMPHYS_BASIC_GEN PARAMS:
+  VDD=1 VSS=0 VTHRESH=0.5
V_V9         N16763641 0 20m
X_U624         N16769550 N16788254 ASYMMETRIC_DELAY PARAMS:
+  RISING_EDGE_DELAY=3u VTHRESH=0.5 FALLING_EDGE_DELAY=3u VDD=1 VSS=0
X_U616         MODE N16761158 N16761170 FPWM COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
R_R1         FB_INT N16761926  200k TC=0,0 
V_V5         N16761170 0 0.8
X_U618         N16761926 N16761940 N16763091 N16769550 COMPHYS_BASIC_GEN
+  PARAMS: VDD=1 VSS=0 VTHRESH=0.5
X_U627         GATE_NMOS GATE_PMOS N16786337 NOR2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U626         SKIP PFM SKIP_PFM_N NAND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
V_V4         N16761158 0 1.2
V_V8         N16763659 0 2m
.ENDS
 
.SUBCKT Pass_Through FB Pass_Through PRECHARGE_ON VIN VOUT  
X_U619         N16774814 PASS_THROUGH_INT N16775115 AND2_BASIC_GEN PARAMS:
+  VDD=1 VSS=0 VTHRESH=500E-3
X_U622         PRECHARGE_ON N16774814 INV_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
V_V5         N16777030 0 582mV
V_V3         N16762684 0 50u
X_U618         N16777030 FB N16762684 N16763662 COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
V_V4         N16776473 0 606mV
X_U615         FB N16776473 N16760966 N16761083 COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
X_U617         N16761083 N16761379 PASS_THROUGH_INT AND2_BASIC_GEN PARAMS:
+  VDD=1 VSS=0 VTHRESH=500E-3
V_V1         N16760966 0 10m
X_U616         VIN VOUT N16771362 N16761379 COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
V_V2         N16771362 0 10m
X_U22         N16775115 N16763662 PASS_THROUGH N16762471 SRLATCHRHP_BASIC_GEN
+  PARAMS: VDD=1 VSS=0 VTHRESH=0.5
.ENDS
 
.SUBCKT OVP OVP VOUT  
V_V2         N16761502 0 0.1
V_V3         N16761602 0 5.7
X_U616         VOUT N16761602 N16761502 OVP COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
.ENDS
 
.SUBCKT Soft_Start FB_INT PRECHARGE_ON SDWN VREF  
X_S69    PRECHARGE_ON 0 SS_TR FB_INT Soft_start_S69 
X_U831         SDWN N16715897 INV_BASIC_GEN PARAMS: VDD=1 VSS=0 VTHRESH=500E-3
X_S68    SDWN 0 SS_TR 0 Soft_start_S68 
E_ABM174         N16734545 0 VALUE {  IF(V(SS_TR) < 0.6, V(SS_TR),0.6)    }
C_C11         VREF 0  10n  TC=0,0 
R_R8         N16734545 VREF  1 TC=0,0 
D_D62         SS_TR N16715923 D_D1 
V_V70         N16715923 0 1
G_ABMII1         N16715923 SS_TR VALUE { IF(V(N16715897) > 0.5,3e-9,0)    }
D_D63         0 SS_TR D_D1 
C_C9         SS_TR 0  5p IC={{SS}*0.6} 
.ENDS
 
.SUBCKT Error_Amp FB ISEN_LDO PFM PRECHARGE_ON REF SDWN VEA  
X_S2    PRECHARGE_ON 0 VEA N16788044 Error_Amp_S2 
R_R6         0 VEA  700MEG TC=0,0 
C_C8         VEA 0  5p  
X_U5         N16784843 VEA D_D
G_ABM2I1         0 VEA VALUE { {LIMIT((V(REF) - V(FB))*7u, -0.5u,0.5u)}    }
V_V8         N16786290 0 295m
X_U6         VEA N16786290 D_D
C_C9         N16782062 0  50p  
E_ABM175         N16788044 0 VALUE { (V(ISEN_LDO) /(0.3*15))    }
X_S1    SDWN 0 VEA 0 Error_Amp_S1 
E_ABM174         N16784843 0 VALUE {  IF(V(PFM) > 0.5, 15m, -95m)    }
R_R4         N16782062 VEA  350k  
.ENDS
 
.SUBCKT Gate_Driver GATE_nMOS GATE_pMOS OVP Pass_Through PRECHARGE PWM PWM_N
+  SDWN SKIP_PFM_N  
C_C10         N16776526 0  1.443n  
C_C7         N16776364 0  1.443n  
X_U630         OVP OVPN INV_BASIC_GEN PARAMS: VDD=1 VSS=0 VTHRESH=500E-3
X_U628         N16794319 N16794600 GATE_NMOS AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U631         LDRV OVPN N16776520 N16794319 AND3_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
R_R7         HDRV N16776526  3  
X_U619         N16776526 N16776520 INV_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
D_D68         LDRV N16776364 D_D1 
X_U620         N16781894 N16782385 INV_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U616         N16776364 N16776358 INV_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U634         SKIP_PFM_N PWM_N N16782385 HDRV AND3_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=500E-3
X_U622         PRECHARGE SDWN N16781894 OR2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U633         SKIP_PFM_N PWM N16802886 LDRV AND3_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U624         PRECHARGE SDWN N16782723 OR2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
D_D69         HDRV N16776526 D_D1 
X_U625         N16782723 N16802886 INV_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U627         PASS_THROUGH N16794600 INV_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
X_U626         N16793571 PASS_THROUGH GATE_PMOS OR2_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=500E-3
R_R5         LDRV N16776364  3  
X_U629         OVPN HDRV N16776358 N16793571 AND3_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
.ENDS
 
.SUBCKT Enable_UVLO EN SDWN VIN VOUT  
E_ABM175         N16761019 0 VALUE {  IF((V(VIN_OK) >0.5 & V(VOUT_OK) > 0.5) ,
+  1.31,  
+ 2m)   }
X_U617         VOUT N16761451 N16761467 VOUT_OK COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
R_R5         EN_INT N16764381  40  
D_D68         N16764381 EN_INT D_D1 
X_U616         VIN N16761003 N16761019 VIN_OK COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
V_V2         N16760737 0 1.2
V_V1         N16760758 0 0.78
V_V4         N16761003 0 1.79
X_U620         N16764381 EN_OK BUF_BASIC_GEN PARAMS: VDD=1 VSS=0 VTHRESH=0.5
V_V5         N16761467 0 10m
X_U618         EN_OK VIN_OK SDWN_N AND2_BASIC_GEN PARAMS: VDD=1 VSS=0
+  VTHRESH=500E-3
C_C7         N16764381 0  1.443u  
X_U615         EN N16760737 N16760758 EN_INT COMPHYS_BASIC_GEN PARAMS: VDD=1
+  VSS=0 VTHRESH=0.5
X_U619         SDWN_N SDWN INV_BASIC_GEN PARAMS: VDD=1 VSS=0 VTHRESH=500E-3
V_V6         N16761451 0 2.19
.ENDS

.subckt TPS61023_schematic_S4 1 2 3 4  
S_S4         3 4 1 2 _S4
RS_S4         1 2 1G
.MODEL         _S4 VSWITCH Roff=100e6 Ron=1m Voff=0.2 Von=0.8
.ends TPS61023_schematic_S4

.subckt TPS61023_schematic_H2 1 2 3 4  
H_H2         3 4 VH_H2 0.3
VH_H2         1 2 0V
.ends TPS61023_schematic_H2

.subckt TPS61023_schematic_S2 1 2 3 4  
S_S2         3 4 1 2 _S2
RS_S2         1 2 1G
.MODEL         _S2 VSWITCH Roff=100MEG Ron=1m Voff=0.2 Von=0.8
.ends TPS61023_schematic_S2

.subckt TPS61023_schematic_S1 1 2 3 4  
S_S1         3 4 1 2 _S1
RS_S1         1 2 1G
.MODEL         _S1 VSWITCH Roff=1e6 Ron=47m Voff=0.2 Von=0.7
.ends TPS61023_schematic_S1

.subckt TPS61023_schematic_F1 1 2 3 4  
F_F1         3 4 VF_F1 1
VF_F1         1 2 0V
.ends TPS61023_schematic_F1

.subckt TPS61023_schematic_H1 1 2 3 4  
H_H1         3 4 VH_H1 0.08
VH_H1         1 2 0V
.ends TPS61023_schematic_H1

.subckt TPS61023_schematic_S3 1 2 3 4  
S_S3         3 4 1 2 _S3
RS_S3         1 2 1G
.MODEL         _S3 VSWITCH Roff=1e6 Ron=68m Voff=0.2 Von=0.7
.ends TPS61023_schematic_S3

.subckt PWM_Control_S2 1 2 3 4  
S_S2         3 4 1 2 _S2
RS_S2         1 2 1G
.MODEL         _S2 VSWITCH Roff=100MEG Ron=20m Voff=0.2 Von=0.8
.ends PWM_Control_S2

.subckt Soft_start_S69 1 2 3 4  
S_S69         3 4 1 2 _S69
RS_S69         1 2 1G
.MODEL         _S69 VSWITCH Roff=100e6 Ron=1m Voff=0.2 Von=0.8
.ends Soft_start_S69

.subckt Soft_start_S68 1 2 3 4  
S_S68         3 4 1 2 _S68
RS_S68         1 2 1G
.MODEL         _S68 VSWITCH Roff=100e9 Ron=1e6 Voff=0.2 Von=0.8
.ends Soft_start_S68

.subckt Error_Amp_S2 1 2 3 4  
S_S2         3 4 1 2 _S2
RS_S2         1 2 1G
.MODEL         _S2 VSWITCH Roff=100MEG Ron=1m Voff=0.2 Von=0.8
.ends Error_Amp_S2

.subckt Error_Amp_S1 1 2 3 4  
S_S1         3 4 1 2 _S1
RS_S1         1 2 1G
.MODEL         _S1 VSWITCH Roff=100MEG Ron=1m Voff=0.2 Von=0.8
.ends Error_Amp_S1

.SUBCKT LDCR IN OUT
+ PARAMS:  L=1u DCR=0.01 IC=0
L	IN 1  {L} IC={IC}
RDCR	1 OUT {DCR}
.ENDS LDCR

.SUBCKT CESR IN OUT
+ PARAMS:  C=100u ESR=0.01 X=1 IC=0
C	IN 1  {C*X} IC={IC}
RESR	1 OUT {ESR/X}
.ENDS CESR

.model D_D1 d
+ is=1e-015
+ n=0.01
+ tt=1e-011

.model MbreakP pmos
+ vto=-0.7
+ kp=10
+ w=4.5e-007
+ l=1e-008
+ lambda=0.12

.subckt d_dnew 1 2
d1 1 2 dd7
.model dd7 d
+ is=1e-015
+ tt=1e-011
+ rs=0.005
+ n=0.01
.ends d_dnew

.SUBCKT INV_BASIC_GEN A  Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 
E_ABMGATE    YINT 0 VALUE {{IF(V(A) > {VTHRESH} , 
+ {VSS},{VDD})}}
RINT YINT Y 1
CINT Y 0 1n
.ENDS INV_BASIC_GEN

.SUBCKT COMP_BASIC_GEN INP INM Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5	
E_ABM Yint 0 VALUE {IF (V(INP) > 
+ V(INM), {VDD},{VSS})}
R1 Yint Y 1
C1 Y 0 1n
.ENDS COMP_BASIC_GEN

.SUBCKT COMPHYS_BASIC_GEN INP INM HYS OUT PARAMS: VDD=1 VSS=0 VTHRESH=0.5	
EIN INP1 INM1 INP INM 1 
EHYS INP1 INP2 VALUE { IF( V(1) > {VTHRESH},-V(HYS),0) }
EOUT OUT 0 VALUE { IF( V(INP2)>V(INM1), {VDD} ,{VSS}) }
R1 OUT 1 1
C1 1 0 5n
RINP1 INP1 0 1K
.ENDS COMPHYS_BASIC_GEN

.SUBCKT AND2_BASIC_GEN A B Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 
E_ABMGATE    YINT 0 VALUE {{IF(V(A) > {VTHRESH}  &  
+ V(B) > {VTHRESH},{VDD},{VSS})}}
RINT YINT Y 1
CINT Y 0 1n
.ENDS AND2_BASIC_GEN

.SUBCKT BUF_BASIC_GEN A  Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 
E_ABMGATE    YINT 0 VALUE {{IF(V(A) > {VTHRESH} , 
+ {VDD},{VSS})}}
RINT YINT Y 1
CINT Y 0 1n
.ENDS BUF_BASIC_GEN

.SUBCKT AND3_BASIC_GEN A B C Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 
E_ABMGATE    YINT 0 VALUE {{IF(V(A) > {VTHRESH}  &  
+ V(B) > {VTHRESH} &
+ V(C) > {VTHRESH},{VDD},{VSS})}}
RINT YINT Y 1
CINT Y 0 1n
.ENDS AND3_BASIC_GEN

.SUBCKT OR2_BASIC_GEN A B Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 
E_ABMGATE    YINT 0 VALUE {{IF(V(A) > {VTHRESH}  |  
+ V(B) > {VTHRESH},{VDD},{VSS})}}
RINT YINT Y 1
CINT Y 0 1n
.ENDS OR2_BASIC_GEN

.subckt d_d 1 2
d1 1 2 dd
.model dd d
+ is=1e-015
+ n=0.01
+ tt=1e-011
.ends d_d

.subckt srlatchrhp_basic_gen s r q qb params: vdd=1 vss=0 vthresh=0.5 
gq 0 qint value = {if(v(r) > {vthresh},-5,if(v(s)>{vthresh},5, 0))}
cqint qint 0 1n
rqint qint 0 1000meg
d_d10 qint my5 d_d1
v1 my5 0 {vdd}
d_d11 myvss qint d_d1
v2 myvss 0 {vss} 
eq qqq 0 qint 0 1
x3 qqq qqqd1 buf_basic_gen params: vdd={vdd} vss={vss} vthresh={vthresh}
rqq qqqd1 q 1
eqb qbr 0 value = {if( v(q) > {vthresh}, {vss},{vdd})}
rqb qbr qb 1 
cdummy1 q 0 1n 
cdummy2 qb 0 1n
.ic v(qint) {vss}
.model d_d1 d
+ is=1e-015
+ tt=1e-011
+ rs=0.05
+ n=0.01
.ends srlatchrhp_basic_gen

.subckt asymmetric_delay inp  out params: rising_edge_delay=1 vthresh=0.5
+  falling_edge_delay=1 vdd=1 vss=0
e_abm3         inp1 0 value { if(v(inp) > {vthresh}, {vdd} , {vss})    }
e_abm1         yin4 0 value { if(v(yin3) > {vthresh}, {vdd} , {vss})    }
e_abm2         yin2 0 value { if(v(yin1) > {vthresh}, {vdd} , {vss})    }
r_rint         inp1 yin1  1  
c_cint         yin1 0  {1.443*rising_edge_delay} 
d_d10         yin1 inp1 d_d1
r_r1         yin4 out  1  
r_rout         yin2 yin3  1  
c_cout         yin3 0 {1.443*falling_edge_delay} 
c_c1         0 out  1n   
d_d11        yin2 yin3 d_d1
.model d_d1 d
+ is=1e-015
+ tt=1e-011
+ rs=0.005
+ n=0.1
.ends asymmetric_delay

.SUBCKT NOR2_BASIC_GEN A B Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 
E_ABMGATE    YINT 0 VALUE {{IF(V(A) > {VTHRESH}  |  
+ V(B) > {VTHRESH},{VSS},{VDD})}}
RINT YINT Y 1
CINT Y 0 1n
.ENDS NOR2_BASIC_GEN

.SUBCKT NAND2_BASIC_GEN A B Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 
E_ABMGATE    YINT 0 VALUE {{IF(V(A) > {VTHRESH}  &  
+ V(B) > {VTHRESH},{VSS},{VDD})}}
RINT YINT Y 1
CINT Y 0 1n
.ENDS NAND2_BASIC_GEN

.SUBCKT INV_DELAY_BASIC_GEN A  Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5 DELAY = 10n 
E_ABMGATE1    YINT1 0 VALUE {{IF(V(A) > {VTHRESH} , 
+ {VDD},{VSS})}}
RINT YINT1 YINT2 1
CINT YINT2 0 {DELAY*1.3}
E_ABMGATE2    YINT3 0 VALUE {{IF(V(YINT2) > {VTHRESH} , 
+ {VSS},{VDD})}}
RINT2 YINT3 Y 1
CINT2 Y 0 1n
.ENDS INV_DELAY_BASIC_GEN

.subckt one_shot in out params:  t=100
s_s1         meas 0 reset2 0 s1
e_abm1         ch 0 value { if( v(in)>0.5 | v(out)>0.5,1,0)    }
r_r2         reset2 reset  0.1  
e_abm3         out 0 value { if( v(meas)<0.5 & v(ch)>0.5,1,0)    }
r_r1         meas ch  {t} 
c_c2         0 reset2  1.4427n  
c_c1         0 meas  1.4427n  
e_abm2         reset 0 value { if(v(ch)<0.5,1,0)    }
.model s1 vswitch
+ roff=1e+009
+ ron=1
+ voff=0.25
+ von=0.75
.ends one_shot

