***********************************************************
*
* PBSS5160T
*
* Nexperia
*
* Low VCEsat PNP (BISS) Transistor
* IC   = 1 A
* VCEO = 60 V 
* hFE  = min. 200 typ. 350 @ 5V/1mA
*
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base
* Package Pin 2: Emitter   
* Package Pin 3: Collector 
*
*
* Extraction date (week/year): 27/2019
* Spicemodel includes temperature dependency
*
**********************************************************
*#
* Please note: Diode D1, Transistor Q2 and Resistor RQ 
* are dedicated to improve modeling of quasi
* saturation area and reverse mode operation
* and do not reflect physical devices.
*
.SUBCKT PBSS5160T B E C
Q1 B E C MAIN 0.881
Q2 11 E C MAIN 0.119
RQ 11 B 16.98
D1 B E DIODE
*
.MODEL MAIN PNP
+ IS = 1.222E-13
+ NF = 0.9536
+ ISE = 8.69E-15
+ NE = 1.272
+ BF = 309.8
+ IKF = 0.6151
+ VAF = 9.213
+ NR = 0.9517
+ ISC = 1.406E-14
+ NC = 1.325
+ BR = 16.64
+ IKR = 7.256
+ VAR = 80
+ RB = 11.5
+ IRB = 0.0008
+ RBM = 2.3
+ RE = 0.07216
+ RC = 0.0612
+ XTB = 1.156
+ EG = 1.11
+ XTI = 2.904
+ CJE = 9.479E-11
+ VJE = 0.7328
+ MJE = 0.3663
+ TF = 1.111E-09
+ XTF = 1.587
+ VTF = 2.697
+ ITF = 0.5379
+ PTF = 0
+ CJC = 3.125E-11
+ VJC = 1
+ MJC = 0.5071
+ XCJC = 1
+ TR = 6.5E-08
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 0.8944
.MODEL DIODE D
+ IS = 8.286E-15
+ N = 0.9998
+ BV = 1000
+ IBV = 0.001
+ RS = 2768
+ CJO = 0
+ VJ = 1
+ M = 0.5
+ FC = 0
+ TT = 0
+ EG = 1.11
+ XTI = 3
.ENDS PBSS5160T
*